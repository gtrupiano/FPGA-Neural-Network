library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.components.all;

entity forward_pass_tb is
end forward_pass_tb;

architecture Behavioral of forward_pass_tb is

signal w1, w2, w3, w4, w5, w6, w7, w8, a1, a2, a3, a4, a5, a6, a7, a8, aout : std_logic_vector(31 downto 0);
signal a_prime : std_logic;

begin

test : Forward_Pass_Neuron_Hidden port map
(
    W1 => w1,
    W2 => w2,
    W3 => w3,
    W4 => w4,
    W5 => w5,
    W6 => w6,
    W7 => w7,
    W8 => w8,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    aout => aout,
    a_prime => a_prime
);

tb : process 
begin
    w1 <= "00000000011110000101000111101011"; --0.47
    w2 <= "00000000111010111000010100011110"; --0.92
    w3 <= "00000000110011110101110000101000"; --0.81
    w4 <= "00000000100011110101110000101000"; --0.56
    w5 <= "00000000110001111010111000010100"; --0.78
    w6 <= "00000000010000000000000000000000"; --0.25
    w7 <= "00000000000101000111101011100001"; --0.08
    w8 <= "00000000011010111000010100011110"; --0.42
    a1 <= "00000000000010100011110101110000"; --0.04
    a2 <= "00000000011000010100011110101110"; --0.38
    a3 <= "00000000111000111101011100001010"; --0.89
    a4 <= "00000000110111000010100011110101"; --0.86
    a5 <= "00000000011101011100001010001111"; --0.46
    a6 <= "00000000100001111010111000010100"; --0.53
    a7 <= "00000000101010001111010111000010"; --0.66
    a8 <= "00000000011000111101011100001010"; --0.39
    wait; --hand calculated output: 2.2788
end process;

end Behavioral;
